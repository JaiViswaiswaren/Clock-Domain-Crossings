`timescale 1ns/1ps
`include "DUAL_FF_SYNC.sv"
`include "WPTR.sv"
`include "RPTR.sv"
`include "ASYNC_FIFO.sv"
